-- soc_system_vip_subsystem.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc_system_vip_subsystem is
	port (
		alt_vip_itc_0_clocked_video_vid_clk          : in  std_logic                      := '0';             --         alt_vip_itc_0_clocked_video.vid_clk
		alt_vip_itc_0_clocked_video_vid_data         : out std_logic_vector(31 downto 0);                     --                                    .vid_data
		alt_vip_itc_0_clocked_video_underflow        : out std_logic;                                         --                                    .underflow
		alt_vip_itc_0_clocked_video_vid_datavalid    : out std_logic;                                         --                                    .vid_datavalid
		alt_vip_itc_0_clocked_video_vid_v_sync       : out std_logic;                                         --                                    .vid_v_sync
		alt_vip_itc_0_clocked_video_vid_h_sync       : out std_logic;                                         --                                    .vid_h_sync
		alt_vip_itc_0_clocked_video_vid_f            : out std_logic;                                         --                                    .vid_f
		alt_vip_itc_0_clocked_video_vid_h            : out std_logic;                                         --                                    .vid_h
		alt_vip_itc_0_clocked_video_vid_v            : out std_logic;                                         --                                    .vid_v
		alt_vip_itc_0_is_clk_rst_clk                 : in  std_logic                      := '0';             --            alt_vip_itc_0_is_clk_rst.clk
		alt_vip_itc_0_is_clk_rst_reset_reset         : in  std_logic                      := '0';             --      alt_vip_itc_0_is_clk_rst_reset.reset
		alt_vip_vfr_hdmi_avalon_master_address       : out std_logic_vector(31 downto 0);                     --      alt_vip_vfr_hdmi_avalon_master.address
		alt_vip_vfr_hdmi_avalon_master_burstcount    : out std_logic_vector(5 downto 0);                      --                                    .burstcount
		alt_vip_vfr_hdmi_avalon_master_readdata      : in  std_logic_vector(127 downto 0) := (others => '0'); --                                    .readdata
		alt_vip_vfr_hdmi_avalon_master_read          : out std_logic;                                         --                                    .read
		alt_vip_vfr_hdmi_avalon_master_readdatavalid : in  std_logic                      := '0';             --                                    .readdatavalid
		alt_vip_vfr_hdmi_avalon_master_waitrequest   : in  std_logic                      := '0';             --                                    .waitrequest
		alt_vip_vfr_hdmi_avalon_slave_address        : in  std_logic_vector(4 downto 0)   := (others => '0'); --       alt_vip_vfr_hdmi_avalon_slave.address
		alt_vip_vfr_hdmi_avalon_slave_write          : in  std_logic                      := '0';             --                                    .write
		alt_vip_vfr_hdmi_avalon_slave_writedata      : in  std_logic_vector(31 downto 0)  := (others => '0'); --                                    .writedata
		alt_vip_vfr_hdmi_avalon_slave_read           : in  std_logic                      := '0';             --                                    .read
		alt_vip_vfr_hdmi_avalon_slave_readdata       : out std_logic_vector(31 downto 0);                     --                                    .readdata
		alt_vip_vfr_hdmi_clock_master_clk            : in  std_logic                      := '0';             --       alt_vip_vfr_hdmi_clock_master.clk
		alt_vip_vfr_hdmi_clock_master_reset_reset    : in  std_logic                      := '0';             -- alt_vip_vfr_hdmi_clock_master_reset.reset
		alt_vip_vfr_hdmi_clock_reset_clk             : in  std_logic                      := '0';             --        alt_vip_vfr_hdmi_clock_reset.clk
		alt_vip_vfr_hdmi_clock_reset_reset_reset     : in  std_logic                      := '0';             --  alt_vip_vfr_hdmi_clock_reset_reset.reset
		alt_vip_vfr_hdmi_interrupt_sender_irq        : out std_logic                                          --   alt_vip_vfr_hdmi_interrupt_sender.irq
	);
end entity soc_system_vip_subsystem;

architecture rtl of soc_system_vip_subsystem is
	component alt_vipitc131_IS2Vid is
		generic (
			NUMBER_OF_COLOUR_PLANES       : integer := 3;
			COLOUR_PLANES_ARE_IN_PARALLEL : integer := 1;
			BPS                           : integer := 8;
			INTERLACED                    : integer := 0;
			H_ACTIVE_PIXELS               : integer := 1920;
			V_ACTIVE_LINES                : integer := 1200;
			ACCEPT_COLOURS_IN_SEQ         : integer := 0;
			FIFO_DEPTH                    : integer := 1920;
			CLOCKS_ARE_SAME               : integer := 0;
			USE_CONTROL                   : integer := 0;
			NO_OF_MODES                   : integer := 1;
			THRESHOLD                     : integer := 1919;
			STD_WIDTH                     : integer := 1;
			GENERATE_SYNC                 : integer := 0;
			USE_EMBEDDED_SYNCS            : integer := 0;
			AP_LINE                       : integer := 0;
			V_BLANK                       : integer := 0;
			H_BLANK                       : integer := 0;
			H_SYNC_LENGTH                 : integer := 44;
			H_FRONT_PORCH                 : integer := 88;
			H_BACK_PORCH                  : integer := 148;
			V_SYNC_LENGTH                 : integer := 5;
			V_FRONT_PORCH                 : integer := 4;
			V_BACK_PORCH                  : integer := 36;
			F_RISING_EDGE                 : integer := 0;
			F_FALLING_EDGE                : integer := 0;
			FIELD0_V_RISING_EDGE          : integer := 0;
			FIELD0_V_BLANK                : integer := 0;
			FIELD0_V_SYNC_LENGTH          : integer := 0;
			FIELD0_V_FRONT_PORCH          : integer := 0;
			FIELD0_V_BACK_PORCH           : integer := 0;
			ANC_LINE                      : integer := 0;
			FIELD0_ANC_LINE               : integer := 0
		);
		port (
			is_clk        : in  std_logic                     := 'X';             -- clk
			rst           : in  std_logic                     := 'X';             -- reset
			is_data       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			is_valid      : in  std_logic                     := 'X';             -- valid
			is_ready      : out std_logic;                                        -- ready
			is_sop        : in  std_logic                     := 'X';             -- startofpacket
			is_eop        : in  std_logic                     := 'X';             -- endofpacket
			vid_clk       : in  std_logic                     := 'X';             -- export
			vid_data      : out std_logic_vector(31 downto 0);                    -- export
			underflow     : out std_logic;                                        -- export
			vid_datavalid : out std_logic;                                        -- export
			vid_v_sync    : out std_logic;                                        -- export
			vid_h_sync    : out std_logic;                                        -- export
			vid_f         : out std_logic;                                        -- export
			vid_h         : out std_logic;                                        -- export
			vid_v         : out std_logic                                         -- export
		);
	end component alt_vipitc131_IS2Vid;

	component alt_vipvfr131_vfr is
		generic (
			BITS_PER_PIXEL_PER_COLOR_PLANE : integer := 8;
			NUMBER_OF_CHANNELS_IN_PARALLEL : integer := 3;
			NUMBER_OF_CHANNELS_IN_SEQUENCE : integer := 1;
			MAX_IMAGE_WIDTH                : integer := 640;
			MAX_IMAGE_HEIGHT               : integer := 480;
			MEM_PORT_WIDTH                 : integer := 256;
			RMASTER_FIFO_DEPTH             : integer := 64;
			RMASTER_BURST_TARGET           : integer := 32;
			CLOCKS_ARE_SEPARATE            : integer := 1
		);
		port (
			clock                : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			master_clock         : in  std_logic                      := 'X';             -- clk
			master_reset         : in  std_logic                      := 'X';             -- reset
			slave_address        : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- address
			slave_write          : in  std_logic                      := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			slave_read           : in  std_logic                      := 'X';             -- read
			slave_readdata       : out std_logic_vector(31 downto 0);                     -- readdata
			slave_irq            : out std_logic;                                         -- irq
			dout_data            : out std_logic_vector(31 downto 0);                     -- data
			dout_valid           : out std_logic;                                         -- valid
			dout_ready           : in  std_logic                      := 'X';             -- ready
			dout_startofpacket   : out std_logic;                                         -- startofpacket
			dout_endofpacket     : out std_logic;                                         -- endofpacket
			master_address       : out std_logic_vector(31 downto 0);                     -- address
			master_burstcount    : out std_logic_vector(5 downto 0);                      -- burstcount
			master_readdata      : in  std_logic_vector(127 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                         -- read
			master_readdatavalid : in  std_logic                      := 'X';             -- readdatavalid
			master_waitrequest   : in  std_logic                      := 'X'              -- waitrequest
		);
	end component alt_vipvfr131_vfr;

	signal alt_vip_vfr_hdmi_avalon_streaming_source_valid         : std_logic;                     -- alt_vip_vfr_hdmi:dout_valid -> alt_vip_itc_0:is_valid
	signal alt_vip_vfr_hdmi_avalon_streaming_source_data          : std_logic_vector(31 downto 0); -- alt_vip_vfr_hdmi:dout_data -> alt_vip_itc_0:is_data
	signal alt_vip_vfr_hdmi_avalon_streaming_source_ready         : std_logic;                     -- alt_vip_itc_0:is_ready -> alt_vip_vfr_hdmi:dout_ready
	signal alt_vip_vfr_hdmi_avalon_streaming_source_startofpacket : std_logic;                     -- alt_vip_vfr_hdmi:dout_startofpacket -> alt_vip_itc_0:is_sop
	signal alt_vip_vfr_hdmi_avalon_streaming_source_endofpacket   : std_logic;                     -- alt_vip_vfr_hdmi:dout_endofpacket -> alt_vip_itc_0:is_eop

begin

	alt_vip_itc_0 : component alt_vipitc131_IS2Vid
		generic map (
			NUMBER_OF_COLOUR_PLANES       => 4,
			COLOUR_PLANES_ARE_IN_PARALLEL => 1,
			BPS                           => 8,
			INTERLACED                    => 0,
			H_ACTIVE_PIXELS               => 1024,
			V_ACTIVE_LINES                => 768,
			ACCEPT_COLOURS_IN_SEQ         => 0,
			FIFO_DEPTH                    => 1920,
			CLOCKS_ARE_SAME               => 0,
			USE_CONTROL                   => 0,
			NO_OF_MODES                   => 1,
			THRESHOLD                     => 1919,
			STD_WIDTH                     => 1,
			GENERATE_SYNC                 => 0,
			USE_EMBEDDED_SYNCS            => 0,
			AP_LINE                       => 0,
			V_BLANK                       => 0,
			H_BLANK                       => 0,
			H_SYNC_LENGTH                 => 136,
			H_FRONT_PORCH                 => 24,
			H_BACK_PORCH                  => 160,
			V_SYNC_LENGTH                 => 6,
			V_FRONT_PORCH                 => 3,
			V_BACK_PORCH                  => 29,
			F_RISING_EDGE                 => 0,
			F_FALLING_EDGE                => 0,
			FIELD0_V_RISING_EDGE          => 0,
			FIELD0_V_BLANK                => 0,
			FIELD0_V_SYNC_LENGTH          => 0,
			FIELD0_V_FRONT_PORCH          => 0,
			FIELD0_V_BACK_PORCH           => 0,
			ANC_LINE                      => 0,
			FIELD0_ANC_LINE               => 0
		)
		port map (
			is_clk        => alt_vip_itc_0_is_clk_rst_clk,                           --       is_clk_rst.clk
			rst           => alt_vip_itc_0_is_clk_rst_reset_reset,                   -- is_clk_rst_reset.reset
			is_data       => alt_vip_vfr_hdmi_avalon_streaming_source_data,          --              din.data
			is_valid      => alt_vip_vfr_hdmi_avalon_streaming_source_valid,         --                 .valid
			is_ready      => alt_vip_vfr_hdmi_avalon_streaming_source_ready,         --                 .ready
			is_sop        => alt_vip_vfr_hdmi_avalon_streaming_source_startofpacket, --                 .startofpacket
			is_eop        => alt_vip_vfr_hdmi_avalon_streaming_source_endofpacket,   --                 .endofpacket
			vid_clk       => alt_vip_itc_0_clocked_video_vid_clk,                    --    clocked_video.export
			vid_data      => alt_vip_itc_0_clocked_video_vid_data,                   --                 .export
			underflow     => alt_vip_itc_0_clocked_video_underflow,                  --                 .export
			vid_datavalid => alt_vip_itc_0_clocked_video_vid_datavalid,              --                 .export
			vid_v_sync    => alt_vip_itc_0_clocked_video_vid_v_sync,                 --                 .export
			vid_h_sync    => alt_vip_itc_0_clocked_video_vid_h_sync,                 --                 .export
			vid_f         => alt_vip_itc_0_clocked_video_vid_f,                      --                 .export
			vid_h         => alt_vip_itc_0_clocked_video_vid_h,                      --                 .export
			vid_v         => alt_vip_itc_0_clocked_video_vid_v                       --                 .export
		);

	alt_vip_vfr_hdmi : component alt_vipvfr131_vfr
		generic map (
			BITS_PER_PIXEL_PER_COLOR_PLANE => 8,
			NUMBER_OF_CHANNELS_IN_PARALLEL => 4,
			NUMBER_OF_CHANNELS_IN_SEQUENCE => 1,
			MAX_IMAGE_WIDTH                => 1024,
			MAX_IMAGE_HEIGHT               => 768,
			MEM_PORT_WIDTH                 => 128,
			RMASTER_FIFO_DEPTH             => 64,
			RMASTER_BURST_TARGET           => 32,
			CLOCKS_ARE_SEPARATE            => 1
		)
		port map (
			clock                => alt_vip_vfr_hdmi_clock_reset_clk,                       --             clock_reset.clk
			reset                => alt_vip_vfr_hdmi_clock_reset_reset_reset,               --       clock_reset_reset.reset
			master_clock         => alt_vip_vfr_hdmi_clock_master_clk,                      --            clock_master.clk
			master_reset         => alt_vip_vfr_hdmi_clock_master_reset_reset,              --      clock_master_reset.reset
			slave_address        => alt_vip_vfr_hdmi_avalon_slave_address,                  --            avalon_slave.address
			slave_write          => alt_vip_vfr_hdmi_avalon_slave_write,                    --                        .write
			slave_writedata      => alt_vip_vfr_hdmi_avalon_slave_writedata,                --                        .writedata
			slave_read           => alt_vip_vfr_hdmi_avalon_slave_read,                     --                        .read
			slave_readdata       => alt_vip_vfr_hdmi_avalon_slave_readdata,                 --                        .readdata
			slave_irq            => alt_vip_vfr_hdmi_interrupt_sender_irq,                  --        interrupt_sender.irq
			dout_data            => alt_vip_vfr_hdmi_avalon_streaming_source_data,          -- avalon_streaming_source.data
			dout_valid           => alt_vip_vfr_hdmi_avalon_streaming_source_valid,         --                        .valid
			dout_ready           => alt_vip_vfr_hdmi_avalon_streaming_source_ready,         --                        .ready
			dout_startofpacket   => alt_vip_vfr_hdmi_avalon_streaming_source_startofpacket, --                        .startofpacket
			dout_endofpacket     => alt_vip_vfr_hdmi_avalon_streaming_source_endofpacket,   --                        .endofpacket
			master_address       => alt_vip_vfr_hdmi_avalon_master_address,                 --           avalon_master.address
			master_burstcount    => alt_vip_vfr_hdmi_avalon_master_burstcount,              --                        .burstcount
			master_readdata      => alt_vip_vfr_hdmi_avalon_master_readdata,                --                        .readdata
			master_read          => alt_vip_vfr_hdmi_avalon_master_read,                    --                        .read
			master_readdatavalid => alt_vip_vfr_hdmi_avalon_master_readdatavalid,           --                        .readdatavalid
			master_waitrequest   => alt_vip_vfr_hdmi_avalon_master_waitrequest              --                        .waitrequest
		);

end architecture rtl; -- of soc_system_vip_subsystem
